
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity I2C_state_tb is
    generic ( 
            DEVICE          : std_logic_vector(7 downto 0) := "01000010"        -- DIRECCI?N DEL DISPOSITIVO 
    );
end I2C_state_tb;

architecture Behavioral of I2C_state_tb is

     constant CLK_PERIOD : time := 8 ns; -- 125 MHz
     signal clk, reset, clr, enable, SDA, NACK, STOP_ACK, OPERA, READ, WRITE, overflow, continue, stop_div : std_logic;
     signal ADDRESS, DATA_IN, DATA_OUT : std_logic_vector(7 downto 0);
     signal div         : std_logic_vector(1 downto 0);

begin

    uut: entity work.I2C_state(Behavioral)
            port map(
                    clk         => clk,
                    reset       => reset,
                    clr         => clr,
                    enable      => enable,
                    SDA         => SDA,
                    ADDRESS     => ADDRESS,
                    DATA_IN     => DATA_IN,
                    DATA_OUT    => DATA_OUT,
                    NACK        => NACK,
                    STOP_ACK    => STOP_ACK,
                    READ        => READ,
                    OPERA       => OPERA,
                    WRITE       => WRITE,
                    overflow    => overflow,
                    div         => div,
                    continue    => continue,
                    stop_div    => stop_div
            );

    clk_stimuli : process
    begin
        clk <= '1';
        wait for CLK_PERIOD/2;
        clk <= '0';
        wait for CLK_PERIOD/2;
    end process;

    uut_stimuli: process
    begin
        -- Se�ales iniciales para causar estado de reset
        reset <= '1';
        OPERA <= '0';
        clr <= '0';
        SDA <= 'Z';
        enable <= '0';
        ADDRESS <= "00000010"; -- Se introducen los bits correspondientes a la direcci�n de memoria del dispositivo
        DATA_IN <= "00000101"; -- Se introducen los bits correspondientes a transmitir en una potencial operaci�n de ESCRITURA
        STOP_ACK <= '0';
        READ <= '0';
        WRITE <= '0';
        overflow <= '0';
        div <= "00";
        wait for 2 us;
    -- Se permite que la parte secuencial trabaje y se introduce el tipo de operaci�n (ESCRITURA)
        WRITE <= '1';
        reset <= '0';
        enable <= '1';
        wait for 2 us;
    -- Se introduce la orden de empezar la operaci�n de ESCRITURA (OPERA funciona a modo de bot�n)
        OPERA <= '1';
        wait for 2 us; -- Se registra la orden (en una se�al intermedia flanco_opera)
        OPERA <= '0';
        
        -- START
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;
                
        -- ESCRITURA DEVICE
        -- 1
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 2
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 3
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 4
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 5
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 6
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 7
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 8
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        -- ACK
        div <= "00";
        wait for 1 us;
        SDA <= '0';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        SDA <= 'Z';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        
        -- ESCRITURA ADDRESS
        -- 1
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 2
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 3
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 4
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';
        wait for 1 us;
        -- 5
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 6
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 7
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 8
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;  
        -- ACK
        div <= "00";
        wait for 1 us;
        SDA <= '0';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        SDA <= 'Z';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;    
         
        -- ESCRITURA DATOS
        -- 1
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 2
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 3
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 4
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';
        wait for 1 us;
        -- 5
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 6
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 7
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 8
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;  
        -- ACK
        div <= "00";
        wait for 1 us;
        SDA <= '0';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        SDA <= 'Z';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        
        -- PRESTOP
        wait for 2 us;
        div <= "00";
        
        -- STOP
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;   
        
        -- IDLE
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;    
        
        -- Se permite que la parte secuencial trabaje y se introduce el tipo de operaci�n (LECTURA)
        WRITE <= '0';
        READ <= '1';
        reset <= '0';
        enable <= '1';
        wait for 2 us;
        -- Se introduce la orden de empezar la operaci�n de LECTURA (OPERA funciona a modo de bot�n)
        OPERA <= '1';
        wait for 2 us; -- Se registra la orden (en una se�al intermedia flanco_opera)
        OPERA <= '0';
            
        -- START
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;   
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;         
        
        -- ESCRITURA DEVICE
        -- 1
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 2
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 3
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 4
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 5
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 6
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 7
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        div <= "00";
        wait for 1 us;
        -- 8
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        -- ACK
        div <= "00";
        wait for 1 us;
        SDA <= '0';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        SDA <= 'Z';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        
        -- ESCRITURA ADDRESS
        -- 1
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 2
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 3
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 4
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';
        wait for 1 us;
        -- 5
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 6
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 7
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 8
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;  
        -- ACK
        div <= "00";
        wait for 1 us;
        SDA <= '0';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        SDA <= 'Z';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;    
         
        -- LECTURA DATOS
        -- 1
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        SDA <= '1';  
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us;
        -- 2
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        SDA <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 3
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        SDA <= '1';  
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 4
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        SDA <= '0';  
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';
        wait for 1 us;
        -- 5
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        SDA <= '1';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 6
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';
        SDA <= '0';    
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        wait for 1 us; 
        -- 7
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        SDA <= '1';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';    
        wait for 1 us;
        -- 8
        div <= "00";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        SDA <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        SDA <= 'Z'; 
        wait for 1 us;  
        -- SENDACK
        div <= "00";
        wait for 1 us;
        --SDA <= '0';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';   
        wait for 1 us;
        div <= "01";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';      
        wait for 1 us;
        div <= "10";
        wait for 1 us;
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';       
        wait for 1 us;
        div <= "11";
        wait for 1 us;
        --SDA <= 'Z';
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0'; 
        
        -- PRESTOP
        wait for 2 us;
        
        -- STOP
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
        wait for 2 us;   
        
        -- IDLE
        overflow <= '1';
        wait for CLK_PERIOD;    
        overflow <= '0';  
                                                                                                                
        wait;
    end process;
end Behavioral;
